magic
tech sky130A
magscale 1 2
timestamp 1729053267
<< viali >>
rect 0 1082 1784 1118
rect 0 36 1784 70
<< metal1 >>
rect -12 1118 1796 1124
rect -12 1082 0 1118
rect 1784 1082 1796 1118
rect -12 1076 1796 1082
rect 166 546 176 598
rect 228 546 238 598
rect 272 550 906 592
rect 950 550 1590 592
rect 1640 546 1650 598
rect 1702 546 1712 598
rect -12 70 1796 76
rect -12 36 0 70
rect 1784 36 1796 70
rect -12 30 1796 36
<< via1 >>
rect 176 546 228 598
rect 1650 546 1702 598
<< metal2 >>
rect 166 598 1712 608
rect 166 546 176 598
rect 228 546 1650 598
rect 1702 546 1712 598
rect 166 538 1712 546
rect 176 536 228 538
rect 1650 536 1702 538
use inverter1  x1
timestamp 1729053267
transform 1 0 54 0 1 616
box -54 -616 369 537
use inverter1  x2
timestamp 1729053267
transform 1 0 733 0 1 616
box -54 -616 369 537
use inverter1  x3
timestamp 1729053267
transform 1 0 1416 0 1 616
box -54 -616 369 537
<< labels >>
flabel viali 10 1106 10 1106 7 FreeSans 800 0 0 0 VDD
port 1 w
flabel viali 16 52 16 52 7 FreeSans 800 0 0 0 GND
port 2 w
flabel via1 1688 576 1688 576 3 FreeSans 800 0 0 0 OUT
port 3 e
<< end >>
