magic
tech sky130A
timestamp 1729047083
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 out
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 gnd
port 2 nsew
<< end >>
